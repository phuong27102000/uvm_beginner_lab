/* ==================================================
 * Filename: top.sv 
 * Date    : 2022-09-24
 * Author  : Nguyen Ha Nhat Phuong
 * Contact : phuong2710@gmail.com
 * ==================================================
 */
module top();
  import uvm_pkg::*;
  import my_pkg::*;

  initial begin
    run_test();
  end
endmodule : top
