/* ==================================================
 * Filename: user_pkg.sv 
 * Date    : 2022-09-24
 * Author  : Nguyen Ha Nhat Phuong
 * Contact : phuong2710@gmail.com
 * ==================================================
 */

package user_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh";
  `include "user_comp.svh";
  `include "user_test.svh";
endpackage : user_pkg
