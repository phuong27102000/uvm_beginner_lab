/*/|==========/=/|====================================/
|*|| Filename |*|| all_components.sv 
|*|| Date     |*|| 2022-12-05
|*|| Author   |*|| Nguyen Ha Nhat Phuong
|*|| Contact  |*|| phuong2710@gmail.com
|_|/==========|_|/===================================*/
`include "components/componentA.sv"
`include "components/componentB.sv"
`include "components/componentC.sv"
`include "components/componentD.sv"
`include "components/componentE.sv"
`include "components/componentF0.sv"
`include "components/componentF1.sv"
`include "components/componentF2.sv"
`include "components/componentG0.sv"
`include "components/componentG1.sv"
`include "components/componentG2.sv"
`include "components/env.sv"
