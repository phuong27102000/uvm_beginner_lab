/*/|==========/=/|====================================/
|*|| Filename |*|| top.sv 
|*|| Date     |*|| 2022-10-09
|*|| Author   |*|| Nguyen Ha Nhat Phuong
|*|| Contact  |*|| phuong2710@gmail.com
|_|/==========|_|/===================================*/

module top;
  import my_pkg ::*;

  initial begin
    run_test("my_test"); 
  end
endmodule: top
