/*/|==========/=/|====================================/
|*|| Filename |*|| test_pkg.sv 
|*|| Date     |*|| 2022-09-29
|*|| Author   |*|| Nguyen Ha Nhat Phuong
|*|| Contact  |*|| phuong2710@gmail.com
|_|/==========|_|/===================================*/

package my_test;
`include "dut_if.sv";
`include "clk_if.sv";
`include "transaction_obj.sv";
`include "generator.sv";
`include "driver.sv";
`include "monitor.sv";
`include "scoreboard.sv";
`include "env.sv";
`include "test.sv"
endpackage : my_test
