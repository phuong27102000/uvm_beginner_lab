/*/|==========/=/|====================================/
|*|| Filename |*|| all_tests.sv 
|*|| Date     |*|| 2022-12-05
|*|| Author   |*|| Nguyen Ha Nhat Phuong
|*|| Contact  |*|| phuong2710@gmail.com
|_|/==========|_|/===================================*/

`include "tests/test.sv";
