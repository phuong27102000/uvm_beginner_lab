/*/|==========/=/|====================================/
|*|| Filename |*|| my_pkg.sv 
|*|| Date     |*|| 2022-09-30
|*|| Author   |*|| Nguyen Ha Nhat Phuong
|*|| Contact  |*|| phuong2710@gmail.com
|_|/==========|_|/===================================*/

package my_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh";
  `include "seq_item.sv";
  `include "sequence.sv";
  `include "driver.sv";
  `include "agent.sv";
  `include "env.sv";
  `include "test.sv";
endpackage : my_pkg
